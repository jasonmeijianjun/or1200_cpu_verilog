library verilog;
use verilog.vl_types.all;
entity or1200_sopc is
    port(
        clk_i           : in     vl_logic;
        rst_i           : in     vl_logic
    );
end or1200_sopc;
