library verilog;
use verilog.vl_types.all;
entity or1200_top is
    generic(
        dw              : integer := 32;
        aw              : integer := 32;
        ppic_ints       : integer := 20;
        boot_adr        : integer := 8388608
    );
    port(
        clk_i           : in     vl_logic;
        rst_i           : in     vl_logic;
        pic_ints_i      : in     vl_logic_vector;
        clmode_i        : in     vl_logic_vector(1 downto 0);
        iwb_clk_i       : in     vl_logic;
        iwb_rst_i       : in     vl_logic;
        iwb_ack_i       : in     vl_logic;
        iwb_err_i       : in     vl_logic;
        iwb_rty_i       : in     vl_logic;
        iwb_dat_i       : in     vl_logic_vector;
        iwb_cyc_o       : out    vl_logic;
        iwb_adr_o       : out    vl_logic_vector;
        iwb_stb_o       : out    vl_logic;
        iwb_we_o        : out    vl_logic;
        iwb_sel_o       : out    vl_logic_vector(3 downto 0);
        iwb_dat_o       : out    vl_logic_vector;
        iwb_cab_o       : out    vl_logic;
        iwb_cti_o       : out    vl_logic_vector(2 downto 0);
        iwb_bte_o       : out    vl_logic_vector(1 downto 0);
        dwb_clk_i       : in     vl_logic;
        dwb_rst_i       : in     vl_logic;
        dwb_ack_i       : in     vl_logic;
        dwb_err_i       : in     vl_logic;
        dwb_rty_i       : in     vl_logic;
        dwb_dat_i       : in     vl_logic_vector;
        dwb_cyc_o       : out    vl_logic;
        dwb_adr_o       : out    vl_logic_vector;
        dwb_stb_o       : out    vl_logic;
        dwb_we_o        : out    vl_logic;
        dwb_sel_o       : out    vl_logic_vector(3 downto 0);
        dwb_dat_o       : out    vl_logic_vector;
        dwb_cab_o       : out    vl_logic;
        dwb_cti_o       : out    vl_logic_vector(2 downto 0);
        dwb_bte_o       : out    vl_logic_vector(1 downto 0);
        dbg_stall_i     : in     vl_logic;
        dbg_ewt_i       : in     vl_logic;
        dbg_lss_o       : out    vl_logic_vector(3 downto 0);
        dbg_is_o        : out    vl_logic_vector(1 downto 0);
        dbg_wp_o        : out    vl_logic_vector(10 downto 0);
        dbg_bp_o        : out    vl_logic;
        dbg_stb_i       : in     vl_logic;
        dbg_we_i        : in     vl_logic;
        dbg_adr_i       : in     vl_logic_vector;
        dbg_dat_i       : in     vl_logic_vector;
        dbg_dat_o       : out    vl_logic_vector;
        dbg_ack_o       : out    vl_logic;
        pm_cpustall_i   : in     vl_logic;
        pm_clksd_o      : out    vl_logic_vector(3 downto 0);
        pm_dc_gate_o    : out    vl_logic;
        pm_ic_gate_o    : out    vl_logic;
        pm_dmmu_gate_o  : out    vl_logic;
        pm_immu_gate_o  : out    vl_logic;
        pm_tt_gate_o    : out    vl_logic;
        pm_cpu_gate_o   : out    vl_logic;
        pm_wakeup_o     : out    vl_logic;
        pm_lvolt_o      : out    vl_logic;
        sig_tick        : out    vl_logic
    );
end or1200_top;
