library verilog;
use verilog.vl_types.all;
entity wb_conmax_slave_if is
    generic(
        pri_sel         : vl_logic_vector(1 downto 0) := (Hi1, Hi0);
        aw              : integer := 32;
        dw              : integer := 32
    );
    port(
        clk_i           : in     vl_logic;
        rst_i           : in     vl_logic;
        conf            : in     vl_logic_vector(15 downto 0);
        wb_data_i       : in     vl_logic_vector;
        wb_data_o       : out    vl_logic_vector;
        wb_addr_o       : out    vl_logic_vector;
        wb_sel_o        : out    vl_logic_vector;
        wb_we_o         : out    vl_logic;
        wb_cyc_o        : out    vl_logic;
        wb_stb_o        : out    vl_logic;
        wb_ack_i        : in     vl_logic;
        wb_err_i        : in     vl_logic;
        wb_rty_i        : in     vl_logic;
        m0_data_i       : in     vl_logic_vector;
        m0_data_o       : out    vl_logic_vector;
        m0_addr_i       : in     vl_logic_vector;
        m0_sel_i        : in     vl_logic_vector;
        m0_we_i         : in     vl_logic;
        m0_cyc_i        : in     vl_logic;
        m0_stb_i        : in     vl_logic;
        m0_ack_o        : out    vl_logic;
        m0_err_o        : out    vl_logic;
        m0_rty_o        : out    vl_logic;
        m1_data_i       : in     vl_logic_vector;
        m1_data_o       : out    vl_logic_vector;
        m1_addr_i       : in     vl_logic_vector;
        m1_sel_i        : in     vl_logic_vector;
        m1_we_i         : in     vl_logic;
        m1_cyc_i        : in     vl_logic;
        m1_stb_i        : in     vl_logic;
        m1_ack_o        : out    vl_logic;
        m1_err_o        : out    vl_logic;
        m1_rty_o        : out    vl_logic;
        m2_data_i       : in     vl_logic_vector;
        m2_data_o       : out    vl_logic_vector;
        m2_addr_i       : in     vl_logic_vector;
        m2_sel_i        : in     vl_logic_vector;
        m2_we_i         : in     vl_logic;
        m2_cyc_i        : in     vl_logic;
        m2_stb_i        : in     vl_logic;
        m2_ack_o        : out    vl_logic;
        m2_err_o        : out    vl_logic;
        m2_rty_o        : out    vl_logic;
        m3_data_i       : in     vl_logic_vector;
        m3_data_o       : out    vl_logic_vector;
        m3_addr_i       : in     vl_logic_vector;
        m3_sel_i        : in     vl_logic_vector;
        m3_we_i         : in     vl_logic;
        m3_cyc_i        : in     vl_logic;
        m3_stb_i        : in     vl_logic;
        m3_ack_o        : out    vl_logic;
        m3_err_o        : out    vl_logic;
        m3_rty_o        : out    vl_logic;
        m4_data_i       : in     vl_logic_vector;
        m4_data_o       : out    vl_logic_vector;
        m4_addr_i       : in     vl_logic_vector;
        m4_sel_i        : in     vl_logic_vector;
        m4_we_i         : in     vl_logic;
        m4_cyc_i        : in     vl_logic;
        m4_stb_i        : in     vl_logic;
        m4_ack_o        : out    vl_logic;
        m4_err_o        : out    vl_logic;
        m4_rty_o        : out    vl_logic;
        m5_data_i       : in     vl_logic_vector;
        m5_data_o       : out    vl_logic_vector;
        m5_addr_i       : in     vl_logic_vector;
        m5_sel_i        : in     vl_logic_vector;
        m5_we_i         : in     vl_logic;
        m5_cyc_i        : in     vl_logic;
        m5_stb_i        : in     vl_logic;
        m5_ack_o        : out    vl_logic;
        m5_err_o        : out    vl_logic;
        m5_rty_o        : out    vl_logic;
        m6_data_i       : in     vl_logic_vector;
        m6_data_o       : out    vl_logic_vector;
        m6_addr_i       : in     vl_logic_vector;
        m6_sel_i        : in     vl_logic_vector;
        m6_we_i         : in     vl_logic;
        m6_cyc_i        : in     vl_logic;
        m6_stb_i        : in     vl_logic;
        m6_ack_o        : out    vl_logic;
        m6_err_o        : out    vl_logic;
        m6_rty_o        : out    vl_logic;
        m7_data_i       : in     vl_logic_vector;
        m7_data_o       : out    vl_logic_vector;
        m7_addr_i       : in     vl_logic_vector;
        m7_sel_i        : in     vl_logic_vector;
        m7_we_i         : in     vl_logic;
        m7_cyc_i        : in     vl_logic;
        m7_stb_i        : in     vl_logic;
        m7_ack_o        : out    vl_logic;
        m7_err_o        : out    vl_logic;
        m7_rty_o        : out    vl_logic
    );
    attribute pri_sel_mti_vect_attrib : integer;
    attribute pri_sel_mti_vect_attrib of pri_sel : constant is 2;
end wb_conmax_slave_if;
