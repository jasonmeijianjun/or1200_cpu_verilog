library verilog;
use verilog.vl_types.all;
entity or1200_except is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic;
        sig_ibuserr     : in     vl_logic;
        sig_dbuserr     : in     vl_logic;
        sig_illegal     : in     vl_logic;
        sig_align       : in     vl_logic;
        sig_range       : in     vl_logic;
        sig_dtlbmiss    : in     vl_logic;
        sig_dmmufault   : in     vl_logic;
        sig_int         : in     vl_logic;
        sig_syscall     : in     vl_logic;
        sig_trap        : in     vl_logic;
        sig_itlbmiss    : in     vl_logic;
        sig_immufault   : in     vl_logic;
        sig_tick        : in     vl_logic;
        ex_branch_taken : in     vl_logic;
        genpc_freeze    : in     vl_logic;
        id_freeze       : in     vl_logic;
        ex_freeze       : in     vl_logic;
        wb_freeze       : in     vl_logic;
        if_stall        : in     vl_logic;
        if_pc           : in     vl_logic_vector(31 downto 0);
        id_pc           : out    vl_logic_vector(31 downto 0);
        ex_pc           : out    vl_logic_vector(31 downto 0);
        wb_pc           : out    vl_logic_vector(31 downto 0);
        id_flushpipe    : in     vl_logic;
        ex_flushpipe    : in     vl_logic;
        extend_flush    : out    vl_logic;
        except_flushpipe: out    vl_logic;
        except_type     : out    vl_logic_vector(3 downto 0);
        except_start    : out    vl_logic;
        except_started  : out    vl_logic;
        except_stop     : out    vl_logic_vector(13 downto 0);
        except_trig     : out    vl_logic_vector(13 downto 0);
        ex_void         : in     vl_logic;
        abort_mvspr     : out    vl_logic;
        branch_op       : in     vl_logic_vector(2 downto 0);
        spr_dat_ppc     : out    vl_logic_vector(31 downto 0);
        spr_dat_npc     : out    vl_logic_vector(31 downto 0);
        datain          : in     vl_logic_vector(31 downto 0);
        du_dsr          : in     vl_logic_vector(13 downto 0);
        epcr_we         : in     vl_logic;
        eear_we         : in     vl_logic;
        esr_we          : in     vl_logic;
        pc_we           : in     vl_logic;
        epcr            : out    vl_logic_vector(31 downto 0);
        eear            : out    vl_logic_vector(31 downto 0);
        du_dmr1         : in     vl_logic_vector(24 downto 0);
        du_hwbkpt       : in     vl_logic;
        du_hwbkpt_ls_r  : in     vl_logic;
        esr             : out    vl_logic_vector(16 downto 0);
        sr_we           : in     vl_logic;
        to_sr           : in     vl_logic_vector(16 downto 0);
        sr              : in     vl_logic_vector(16 downto 0);
        lsu_addr        : in     vl_logic_vector(31 downto 0);
        abort_ex        : out    vl_logic;
        icpu_ack_i      : in     vl_logic;
        icpu_err_i      : in     vl_logic;
        dcpu_ack_i      : in     vl_logic;
        dcpu_err_i      : in     vl_logic;
        sig_fp          : in     vl_logic;
        fpcsr_fpee      : in     vl_logic
    );
end or1200_except;
