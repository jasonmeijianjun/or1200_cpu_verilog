library verilog;
use verilog.vl_types.all;
entity wb_conmax_master_if is
    generic(
        dw              : integer := 32;
        aw              : integer := 32
    );
    port(
        clk_i           : in     vl_logic;
        rst_i           : in     vl_logic;
        wb_data_i       : in     vl_logic_vector;
        wb_data_o       : out    vl_logic_vector;
        wb_addr_i       : in     vl_logic_vector;
        wb_sel_i        : in     vl_logic_vector;
        wb_we_i         : in     vl_logic;
        wb_cyc_i        : in     vl_logic;
        wb_stb_i        : in     vl_logic;
        wb_ack_o        : out    vl_logic;
        wb_err_o        : out    vl_logic;
        wb_rty_o        : out    vl_logic;
        s0_data_i       : in     vl_logic_vector;
        s0_data_o       : out    vl_logic_vector;
        s0_addr_o       : out    vl_logic_vector;
        s0_sel_o        : out    vl_logic_vector;
        s0_we_o         : out    vl_logic;
        s0_cyc_o        : out    vl_logic;
        s0_stb_o        : out    vl_logic;
        s0_ack_i        : in     vl_logic;
        s0_err_i        : in     vl_logic;
        s0_rty_i        : in     vl_logic;
        s1_data_i       : in     vl_logic_vector;
        s1_data_o       : out    vl_logic_vector;
        s1_addr_o       : out    vl_logic_vector;
        s1_sel_o        : out    vl_logic_vector;
        s1_we_o         : out    vl_logic;
        s1_cyc_o        : out    vl_logic;
        s1_stb_o        : out    vl_logic;
        s1_ack_i        : in     vl_logic;
        s1_err_i        : in     vl_logic;
        s1_rty_i        : in     vl_logic;
        s2_data_i       : in     vl_logic_vector;
        s2_data_o       : out    vl_logic_vector;
        s2_addr_o       : out    vl_logic_vector;
        s2_sel_o        : out    vl_logic_vector;
        s2_we_o         : out    vl_logic;
        s2_cyc_o        : out    vl_logic;
        s2_stb_o        : out    vl_logic;
        s2_ack_i        : in     vl_logic;
        s2_err_i        : in     vl_logic;
        s2_rty_i        : in     vl_logic;
        s3_data_i       : in     vl_logic_vector;
        s3_data_o       : out    vl_logic_vector;
        s3_addr_o       : out    vl_logic_vector;
        s3_sel_o        : out    vl_logic_vector;
        s3_we_o         : out    vl_logic;
        s3_cyc_o        : out    vl_logic;
        s3_stb_o        : out    vl_logic;
        s3_ack_i        : in     vl_logic;
        s3_err_i        : in     vl_logic;
        s3_rty_i        : in     vl_logic;
        s4_data_i       : in     vl_logic_vector;
        s4_data_o       : out    vl_logic_vector;
        s4_addr_o       : out    vl_logic_vector;
        s4_sel_o        : out    vl_logic_vector;
        s4_we_o         : out    vl_logic;
        s4_cyc_o        : out    vl_logic;
        s4_stb_o        : out    vl_logic;
        s4_ack_i        : in     vl_logic;
        s4_err_i        : in     vl_logic;
        s4_rty_i        : in     vl_logic;
        s5_data_i       : in     vl_logic_vector;
        s5_data_o       : out    vl_logic_vector;
        s5_addr_o       : out    vl_logic_vector;
        s5_sel_o        : out    vl_logic_vector;
        s5_we_o         : out    vl_logic;
        s5_cyc_o        : out    vl_logic;
        s5_stb_o        : out    vl_logic;
        s5_ack_i        : in     vl_logic;
        s5_err_i        : in     vl_logic;
        s5_rty_i        : in     vl_logic;
        s6_data_i       : in     vl_logic_vector;
        s6_data_o       : out    vl_logic_vector;
        s6_addr_o       : out    vl_logic_vector;
        s6_sel_o        : out    vl_logic_vector;
        s6_we_o         : out    vl_logic;
        s6_cyc_o        : out    vl_logic;
        s6_stb_o        : out    vl_logic;
        s6_ack_i        : in     vl_logic;
        s6_err_i        : in     vl_logic;
        s6_rty_i        : in     vl_logic;
        s7_data_i       : in     vl_logic_vector;
        s7_data_o       : out    vl_logic_vector;
        s7_addr_o       : out    vl_logic_vector;
        s7_sel_o        : out    vl_logic_vector;
        s7_we_o         : out    vl_logic;
        s7_cyc_o        : out    vl_logic;
        s7_stb_o        : out    vl_logic;
        s7_ack_i        : in     vl_logic;
        s7_err_i        : in     vl_logic;
        s7_rty_i        : in     vl_logic;
        s8_data_i       : in     vl_logic_vector;
        s8_data_o       : out    vl_logic_vector;
        s8_addr_o       : out    vl_logic_vector;
        s8_sel_o        : out    vl_logic_vector;
        s8_we_o         : out    vl_logic;
        s8_cyc_o        : out    vl_logic;
        s8_stb_o        : out    vl_logic;
        s8_ack_i        : in     vl_logic;
        s8_err_i        : in     vl_logic;
        s8_rty_i        : in     vl_logic;
        s9_data_i       : in     vl_logic_vector;
        s9_data_o       : out    vl_logic_vector;
        s9_addr_o       : out    vl_logic_vector;
        s9_sel_o        : out    vl_logic_vector;
        s9_we_o         : out    vl_logic;
        s9_cyc_o        : out    vl_logic;
        s9_stb_o        : out    vl_logic;
        s9_ack_i        : in     vl_logic;
        s9_err_i        : in     vl_logic;
        s9_rty_i        : in     vl_logic;
        s10_data_i      : in     vl_logic_vector;
        s10_data_o      : out    vl_logic_vector;
        s10_addr_o      : out    vl_logic_vector;
        s10_sel_o       : out    vl_logic_vector;
        s10_we_o        : out    vl_logic;
        s10_cyc_o       : out    vl_logic;
        s10_stb_o       : out    vl_logic;
        s10_ack_i       : in     vl_logic;
        s10_err_i       : in     vl_logic;
        s10_rty_i       : in     vl_logic;
        s11_data_i      : in     vl_logic_vector;
        s11_data_o      : out    vl_logic_vector;
        s11_addr_o      : out    vl_logic_vector;
        s11_sel_o       : out    vl_logic_vector;
        s11_we_o        : out    vl_logic;
        s11_cyc_o       : out    vl_logic;
        s11_stb_o       : out    vl_logic;
        s11_ack_i       : in     vl_logic;
        s11_err_i       : in     vl_logic;
        s11_rty_i       : in     vl_logic;
        s12_data_i      : in     vl_logic_vector;
        s12_data_o      : out    vl_logic_vector;
        s12_addr_o      : out    vl_logic_vector;
        s12_sel_o       : out    vl_logic_vector;
        s12_we_o        : out    vl_logic;
        s12_cyc_o       : out    vl_logic;
        s12_stb_o       : out    vl_logic;
        s12_ack_i       : in     vl_logic;
        s12_err_i       : in     vl_logic;
        s12_rty_i       : in     vl_logic;
        s13_data_i      : in     vl_logic_vector;
        s13_data_o      : out    vl_logic_vector;
        s13_addr_o      : out    vl_logic_vector;
        s13_sel_o       : out    vl_logic_vector;
        s13_we_o        : out    vl_logic;
        s13_cyc_o       : out    vl_logic;
        s13_stb_o       : out    vl_logic;
        s13_ack_i       : in     vl_logic;
        s13_err_i       : in     vl_logic;
        s13_rty_i       : in     vl_logic;
        s14_data_i      : in     vl_logic_vector;
        s14_data_o      : out    vl_logic_vector;
        s14_addr_o      : out    vl_logic_vector;
        s14_sel_o       : out    vl_logic_vector;
        s14_we_o        : out    vl_logic;
        s14_cyc_o       : out    vl_logic;
        s14_stb_o       : out    vl_logic;
        s14_ack_i       : in     vl_logic;
        s14_err_i       : in     vl_logic;
        s14_rty_i       : in     vl_logic;
        s15_data_i      : in     vl_logic_vector;
        s15_data_o      : out    vl_logic_vector;
        s15_addr_o      : out    vl_logic_vector;
        s15_sel_o       : out    vl_logic_vector;
        s15_we_o        : out    vl_logic;
        s15_cyc_o       : out    vl_logic;
        s15_stb_o       : out    vl_logic;
        s15_ack_i       : in     vl_logic;
        s15_err_i       : in     vl_logic;
        s15_rty_i       : in     vl_logic
    );
end wb_conmax_master_if;
