library verilog;
use verilog.vl_types.all;
entity or1200_sopc_tb is
end or1200_sopc_tb;
